
module SP_unit (
	source,
	probe,
	source_clk);	

	output	[0:0]	source;
	input	[9:0]	probe;
	input		source_clk;
endmodule
