
module SP_unit (
	source,
	source_clk);	

	output	[8:0]	source;
	input		source_clk;
endmodule
