`timescale 1 ns / 1 ns
module lab_PD3_top (
	input bit clk,
	input bit reset,
	output bit [7:0] ledA,
	output bit [31:0] ledB
);
lab_PD3 lab3_1_inst (
	.clk_clk       (clk),   
	.reset_reset_n (reset), 
	.dout_a_export (ledA),  
	.dout_b_export (ledB)   
);
endmodule
