
module lab_PD2 (
	clk_clk,
	reset_reset_n,
	dout_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	dout_export;
endmodule
