module mult_LP_V1 #(
  parameter W = 4
) (
  input                clk,         // Входной тактовый сигнал
  input      [  W-1:0] dA,          // Входной операнд A
  input      [  W-1:0] dB,          // Входной операнд B
  output reg [2*W-1:0] a_mult_b     // Выход, хранящий результат умножения
);

  reg [2*W-1:0] dSUM[0:W];           // Массив для хранения промежуточных результатов суммы
  reg [  W-1:0] A   [0:W];           // Массив для хранения промежуточных значений операнда A
  reg [  W-1:0] B   [0:W];           // Массив для хранения промежуточных значений операнда B

  // Начальные значения для массивов и результата
  initial begin
    for (int i = 0; i <= W; i++) begin
      dSUM[i] <= 1'b0;
      A[i]    <= 1'b0;
      B[i]    <= 1'b0;
    end
    a_mult_b <= 1'b0;
  end

  // На каждом положительном фронте тактового сигнала, присваиваем значения dA и dB соответственно в A[0] и B[0]
  always @(posedge clk) begin
    A[0] <= dA;
    B[0] <= dB;
  end

  genvar i;
  generate
    // Используем генерацию кода для создания параллельных блоков (генераторов) для каждого бита входного операнда
    for (i = 0; i < W; i++) begin : generator
      // На каждом положительном фронте тактового сигнала, обновляем промежуточные значения dSUM, A и B
      always @(posedge clk) begin
        dSUM[i+1] <= (dSUM[i] << 1'b1) + (B[i][W-i-1] ? A[i] : 1'b0);
        A[i+1]    <= A[i];
        B[i+1]    <= B[i];
      end
    end
  endgenerate

  // На каждом положительном фронте тактового сигнала, присваиваем значение dSUM[W] регистру a_mult_b
  always @(posedge clk) a_mult_b <= dSUM[W];

endmodule
