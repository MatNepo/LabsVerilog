
module sp_unit (
	source,
	probe,
	source_clk);	

	output	[18:0]	source;
	input	[7:0]	probe;
	input		source_clk;
endmodule
