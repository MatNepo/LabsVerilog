
module SP (
	source,
	source_clk);	

	output	[0:0]	source;
	input		source_clk;
endmodule
