// lab_PD1_sys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module lab_PD1_sys (
		output wire [31:0] alu0_out_data,   //  alu0_out.data
		input  wire        alu0_out_ready,  //          .ready
		output wire        alu0_out_valid,  //          .valid
		output wire [31:0] alu1_out_data,   //  alu1_out.data
		input  wire        alu1_out_ready,  //          .ready
		output wire        alu1_out_valid,  //          .valid
		input  wire        clk_clk,         //       clk.clk
		output wire        delay_out_valid, // delay_out.valid
		output wire [31:0] delay_out_data,  //          .data
		input  wire        reset_reset_n    //     reset.reset_n
	);

	wire         mm_stream_source_out0_valid;                       // MM_Stream_source:aso_out0_valid -> st_splitter:in0_valid
	wire  [31:0] mm_stream_source_out0_data;                        // MM_Stream_source:aso_out0_data -> st_splitter:in0_data
	wire         mm_stream_source_out0_ready;                       // st_splitter:in0_ready -> MM_Stream_source:aso_out0_ready
	wire         st_splitter_out0_valid;                            // st_splitter:out0_valid -> ST_ALU_1:asi_in1_valid
	wire  [31:0] st_splitter_out0_data;                             // st_splitter:out0_data -> ST_ALU_1:asi_in1_data
	wire         st_splitter_out0_ready;                            // ST_ALU_1:asi_in1_ready -> st_splitter:out0_ready
	wire         st_splitter_out1_valid;                            // st_splitter:out1_valid -> ST_ALU_1:asi_in0_valid
	wire  [31:0] st_splitter_out1_data;                             // st_splitter:out1_data -> ST_ALU_1:asi_in0_data
	wire         st_splitter_out1_ready;                            // ST_ALU_1:asi_in0_ready -> st_splitter:out1_ready
	wire         st_splitter_out2_valid;                            // st_splitter:out2_valid -> ST_ALU_0:asi_in1_valid
	wire  [31:0] st_splitter_out2_data;                             // st_splitter:out2_data -> ST_ALU_0:asi_in1_data
	wire         st_splitter_out2_ready;                            // ST_ALU_0:asi_in1_ready -> st_splitter:out2_ready
	wire         st_splitter_out3_valid;                            // st_splitter:out3_valid -> ST_ALU_0:asi_in0_valid
	wire  [31:0] st_splitter_out3_data;                             // st_splitter:out3_data -> ST_ALU_0:asi_in0_data
	wire         st_splitter_out3_ready;                            // ST_ALU_0:asi_in0_ready -> st_splitter:out3_ready
	wire         my_masterb_m0_waitrequest;                         // mm_interconnect_0:my_masterB_m0_waitrequest -> my_masterB:avm_m0_waitrequest
	wire  [31:0] my_masterb_m0_address;                             // my_masterB:avm_m0_address -> mm_interconnect_0:my_masterB_m0_address
	wire         my_masterb_m0_write;                               // my_masterB:avm_m0_write -> mm_interconnect_0:my_masterB_m0_write
	wire  [31:0] my_masterb_m0_writedata;                           // my_masterB:avm_m0_writedata -> mm_interconnect_0:my_masterB_m0_writedata
	wire         mm_interconnect_0_st_alu_0_s0_waitrequest;         // ST_ALU_0:avs_s0_waitrequest -> mm_interconnect_0:ST_ALU_0_s0_waitrequest
	wire         mm_interconnect_0_st_alu_0_s0_write;               // mm_interconnect_0:ST_ALU_0_s0_write -> ST_ALU_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_st_alu_0_s0_writedata;           // mm_interconnect_0:ST_ALU_0_s0_writedata -> ST_ALU_0:avs_s0_writedata
	wire         mm_interconnect_0_st_alu_1_s0_waitrequest;         // ST_ALU_1:avs_s0_waitrequest -> mm_interconnect_0:ST_ALU_1_s0_waitrequest
	wire         mm_interconnect_0_st_alu_1_s0_write;               // mm_interconnect_0:ST_ALU_1_s0_write -> ST_ALU_1:avs_s0_write
	wire  [31:0] mm_interconnect_0_st_alu_1_s0_writedata;           // mm_interconnect_0:ST_ALU_1_s0_writedata -> ST_ALU_1:avs_s0_writedata
	wire         my_mastera_m0_waitrequest;                         // mm_interconnect_1:my_masterA_m0_waitrequest -> my_masterA:avm_m0_waitrequest
	wire  [31:0] my_mastera_m0_address;                             // my_masterA:avm_m0_address -> mm_interconnect_1:my_masterA_m0_address
	wire         my_mastera_m0_write;                               // my_masterA:avm_m0_write -> mm_interconnect_1:my_masterA_m0_write
	wire  [31:0] my_mastera_m0_writedata;                           // my_masterA:avm_m0_writedata -> mm_interconnect_1:my_masterA_m0_writedata
	wire         mm_interconnect_1_mm_stream_source_s0_waitrequest; // MM_Stream_source:avs_s0_waitrequest -> mm_interconnect_1:MM_Stream_source_s0_waitrequest
	wire         mm_interconnect_1_mm_stream_source_s0_write;       // mm_interconnect_1:MM_Stream_source_s0_write -> MM_Stream_source:avs_s0_write
	wire  [31:0] mm_interconnect_1_mm_stream_source_s0_writedata;   // mm_interconnect_1:MM_Stream_source_s0_writedata -> MM_Stream_source:avs_s0_writedata
	wire         st_splitter_out4_valid;                            // st_splitter:out4_valid -> avalon_st_adapter:in_0_valid
	wire  [31:0] st_splitter_out4_data;                             // st_splitter:out4_data -> avalon_st_adapter:in_0_data
	wire         st_splitter_out4_ready;                            // avalon_st_adapter:in_0_ready -> st_splitter:out4_ready
	wire         avalon_st_adapter_out_0_valid;                     // avalon_st_adapter:out_0_valid -> st_delay:in0_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                      // avalon_st_adapter:out_0_data -> st_delay:in0_data

	MM_Stream_source mm_stream_source (
		.csi_clk            (clk_clk),                                           // clock.clk
		.rsi_reset          (~reset_reset_n),                                    // reset.reset
		.aso_out0_data      (mm_stream_source_out0_data),                        //  out0.data
		.aso_out0_ready     (mm_stream_source_out0_ready),                       //      .ready
		.aso_out0_valid     (mm_stream_source_out0_valid),                       //      .valid
		.avs_s0_writedata   (mm_interconnect_1_mm_stream_source_s0_writedata),   //    s0.writedata
		.avs_s0_write       (mm_interconnect_1_mm_stream_source_s0_write),       //      .write
		.avs_s0_waitrequest (mm_interconnect_1_mm_stream_source_s0_waitrequest)  //      .waitrequest
	);

	ST_ALU st_alu_0 (
		.csi_clk            (clk_clk),                                   // clock.clk
		.rsi_reset          (~reset_reset_n),                            // reset.reset
		.asi_in0_data       (st_splitter_out3_data),                     //   in0.data
		.asi_in0_valid      (st_splitter_out3_valid),                    //      .valid
		.asi_in0_ready      (st_splitter_out3_ready),                    //      .ready
		.asi_in1_data       (st_splitter_out2_data),                     //   in1.data
		.asi_in1_valid      (st_splitter_out2_valid),                    //      .valid
		.asi_in1_ready      (st_splitter_out2_ready),                    //      .ready
		.aso_out0_data      (alu0_out_data),                             //  out0.data
		.aso_out0_ready     (alu0_out_ready),                            //      .ready
		.aso_out0_valid     (alu0_out_valid),                            //      .valid
		.avs_s0_writedata   (mm_interconnect_0_st_alu_0_s0_writedata),   //    s0.writedata
		.avs_s0_write       (mm_interconnect_0_st_alu_0_s0_write),       //      .write
		.avs_s0_waitrequest (mm_interconnect_0_st_alu_0_s0_waitrequest)  //      .waitrequest
	);

	ST_ALU st_alu_1 (
		.csi_clk            (clk_clk),                                   // clock.clk
		.rsi_reset          (~reset_reset_n),                            // reset.reset
		.asi_in0_data       (st_splitter_out1_data),                     //   in0.data
		.asi_in0_valid      (st_splitter_out1_valid),                    //      .valid
		.asi_in0_ready      (st_splitter_out1_ready),                    //      .ready
		.asi_in1_data       (st_splitter_out0_data),                     //   in1.data
		.asi_in1_valid      (st_splitter_out0_valid),                    //      .valid
		.asi_in1_ready      (st_splitter_out0_ready),                    //      .ready
		.aso_out0_data      (alu1_out_data),                             //  out0.data
		.aso_out0_ready     (alu1_out_ready),                            //      .ready
		.aso_out0_valid     (alu1_out_valid),                            //      .valid
		.avs_s0_writedata   (mm_interconnect_0_st_alu_1_s0_writedata),   //    s0.writedata
		.avs_s0_write       (mm_interconnect_0_st_alu_1_s0_write),       //      .write
		.avs_s0_waitrequest (mm_interconnect_0_st_alu_1_s0_waitrequest)  //      .waitrequest
	);

	my_masterA #(
		.address (0),
		.data    (100)
	) my_mastera (
		.csi_clk            (clk_clk),                   // clock.clk
		.rsi_reset          (~reset_reset_n),            // reset.reset
		.avm_m0_address     (my_mastera_m0_address),     //    m0.address
		.avm_m0_write       (my_mastera_m0_write),       //      .write
		.avm_m0_writedata   (my_mastera_m0_writedata),   //      .writedata
		.avm_m0_waitrequest (my_mastera_m0_waitrequest)  //      .waitrequest
	);

	my_masterB #(
		.address_1 (0),
		.data_1    (111),
		.address_2 (4),
		.data_2    (222)
	) my_masterb (
		.csi_clk            (clk_clk),                   // clock.clk
		.rsi_reset          (~reset_reset_n),            // reset.reset
		.avm_m0_address     (my_masterb_m0_address),     //    m0.address
		.avm_m0_write       (my_masterb_m0_write),       //      .write
		.avm_m0_writedata   (my_masterb_m0_writedata),   //      .writedata
		.avm_m0_waitrequest (my_masterb_m0_waitrequest)  //      .waitrequest
	);

	altera_avalon_st_delay #(
		.NUMBER_OF_DELAY_CLOCKS (1),
		.DATA_WIDTH             (32),
		.BITS_PER_SYMBOL        (8),
		.USE_PACKETS            (0),
		.USE_CHANNEL            (0),
		.CHANNEL_WIDTH          (1),
		.USE_ERROR              (0),
		.ERROR_WIDTH            (1)
	) st_delay (
		.in0_valid          (avalon_st_adapter_out_0_valid), //        in.valid
		.in0_data           (avalon_st_adapter_out_0_data),  //          .data
		.out0_valid         (delay_out_valid),               //       out.valid
		.out0_data          (delay_out_data),                //          .data
		.clk                (clk_clk),                       //       clk.clk
		.reset_n            (reset_reset_n),                 // clk_reset.reset_n
		.in0_startofpacket  (1'b0),                          // (terminated)
		.in0_endofpacket    (1'b0),                          // (terminated)
		.out0_startofpacket (),                              // (terminated)
		.out0_endofpacket   (),                              // (terminated)
		.in0_empty          (1'b0),                          // (terminated)
		.out0_empty         (),                              // (terminated)
		.in0_channel        (1'b0),                          // (terminated)
		.out0_channel       (),                              // (terminated)
		.in0_error          (1'b0),                          // (terminated)
		.out0_error         ()                               // (terminated)
	);

	altera_avalon_st_splitter #(
		.NUMBER_OF_OUTPUTS (5),
		.QUALIFY_VALID_OUT (1),
		.USE_PACKETS       (0),
		.DATA_WIDTH        (32),
		.CHANNEL_WIDTH     (1),
		.ERROR_WIDTH       (1),
		.BITS_PER_SYMBOL   (8),
		.EMPTY_WIDTH       (2)
	) st_splitter (
		.clk                 (clk_clk),                     //   clk.clk
		.reset               (~reset_reset_n),              // reset.reset
		.in0_ready           (mm_stream_source_out0_ready), //    in.ready
		.in0_valid           (mm_stream_source_out0_valid), //      .valid
		.in0_data            (mm_stream_source_out0_data),  //      .data
		.out0_ready          (st_splitter_out0_ready),      //  out0.ready
		.out0_valid          (st_splitter_out0_valid),      //      .valid
		.out0_data           (st_splitter_out0_data),       //      .data
		.out1_ready          (st_splitter_out1_ready),      //  out1.ready
		.out1_valid          (st_splitter_out1_valid),      //      .valid
		.out1_data           (st_splitter_out1_data),       //      .data
		.out2_ready          (st_splitter_out2_ready),      //  out2.ready
		.out2_valid          (st_splitter_out2_valid),      //      .valid
		.out2_data           (st_splitter_out2_data),       //      .data
		.out3_ready          (st_splitter_out3_ready),      //  out3.ready
		.out3_valid          (st_splitter_out3_valid),      //      .valid
		.out3_data           (st_splitter_out3_data),       //      .data
		.out4_ready          (st_splitter_out4_ready),      //  out4.ready
		.out4_valid          (st_splitter_out4_valid),      //      .valid
		.out4_data           (st_splitter_out4_data),       //      .data
		.in0_startofpacket   (1'b0),                        // (terminated)
		.in0_endofpacket     (1'b0),                        // (terminated)
		.in0_empty           (2'b00),                       // (terminated)
		.in0_channel         (1'b0),                        // (terminated)
		.in0_error           (1'b0),                        // (terminated)
		.out0_startofpacket  (),                            // (terminated)
		.out0_endofpacket    (),                            // (terminated)
		.out0_empty          (),                            // (terminated)
		.out0_channel        (),                            // (terminated)
		.out0_error          (),                            // (terminated)
		.out1_startofpacket  (),                            // (terminated)
		.out1_endofpacket    (),                            // (terminated)
		.out1_empty          (),                            // (terminated)
		.out1_channel        (),                            // (terminated)
		.out1_error          (),                            // (terminated)
		.out2_startofpacket  (),                            // (terminated)
		.out2_endofpacket    (),                            // (terminated)
		.out2_empty          (),                            // (terminated)
		.out2_channel        (),                            // (terminated)
		.out2_error          (),                            // (terminated)
		.out3_startofpacket  (),                            // (terminated)
		.out3_endofpacket    (),                            // (terminated)
		.out3_empty          (),                            // (terminated)
		.out3_channel        (),                            // (terminated)
		.out3_error          (),                            // (terminated)
		.out4_startofpacket  (),                            // (terminated)
		.out4_endofpacket    (),                            // (terminated)
		.out4_empty          (),                            // (terminated)
		.out4_channel        (),                            // (terminated)
		.out4_error          (),                            // (terminated)
		.out5_ready          (1'b1),                        // (terminated)
		.out5_valid          (),                            // (terminated)
		.out5_startofpacket  (),                            // (terminated)
		.out5_endofpacket    (),                            // (terminated)
		.out5_empty          (),                            // (terminated)
		.out5_channel        (),                            // (terminated)
		.out5_error          (),                            // (terminated)
		.out5_data           (),                            // (terminated)
		.out6_ready          (1'b1),                        // (terminated)
		.out6_valid          (),                            // (terminated)
		.out6_startofpacket  (),                            // (terminated)
		.out6_endofpacket    (),                            // (terminated)
		.out6_empty          (),                            // (terminated)
		.out6_channel        (),                            // (terminated)
		.out6_error          (),                            // (terminated)
		.out6_data           (),                            // (terminated)
		.out7_ready          (1'b1),                        // (terminated)
		.out7_valid          (),                            // (terminated)
		.out7_startofpacket  (),                            // (terminated)
		.out7_endofpacket    (),                            // (terminated)
		.out7_empty          (),                            // (terminated)
		.out7_channel        (),                            // (terminated)
		.out7_error          (),                            // (terminated)
		.out7_data           (),                            // (terminated)
		.out8_ready          (1'b1),                        // (terminated)
		.out8_valid          (),                            // (terminated)
		.out8_startofpacket  (),                            // (terminated)
		.out8_endofpacket    (),                            // (terminated)
		.out8_empty          (),                            // (terminated)
		.out8_channel        (),                            // (terminated)
		.out8_error          (),                            // (terminated)
		.out8_data           (),                            // (terminated)
		.out9_ready          (1'b1),                        // (terminated)
		.out9_valid          (),                            // (terminated)
		.out9_startofpacket  (),                            // (terminated)
		.out9_endofpacket    (),                            // (terminated)
		.out9_empty          (),                            // (terminated)
		.out9_channel        (),                            // (terminated)
		.out9_error          (),                            // (terminated)
		.out9_data           (),                            // (terminated)
		.out10_ready         (1'b1),                        // (terminated)
		.out10_valid         (),                            // (terminated)
		.out10_startofpacket (),                            // (terminated)
		.out10_endofpacket   (),                            // (terminated)
		.out10_empty         (),                            // (terminated)
		.out10_channel       (),                            // (terminated)
		.out10_error         (),                            // (terminated)
		.out10_data          (),                            // (terminated)
		.out11_ready         (1'b1),                        // (terminated)
		.out11_valid         (),                            // (terminated)
		.out11_startofpacket (),                            // (terminated)
		.out11_endofpacket   (),                            // (terminated)
		.out11_empty         (),                            // (terminated)
		.out11_channel       (),                            // (terminated)
		.out11_error         (),                            // (terminated)
		.out11_data          (),                            // (terminated)
		.out12_ready         (1'b1),                        // (terminated)
		.out12_valid         (),                            // (terminated)
		.out12_startofpacket (),                            // (terminated)
		.out12_endofpacket   (),                            // (terminated)
		.out12_empty         (),                            // (terminated)
		.out12_channel       (),                            // (terminated)
		.out12_error         (),                            // (terminated)
		.out12_data          (),                            // (terminated)
		.out13_ready         (1'b1),                        // (terminated)
		.out13_valid         (),                            // (terminated)
		.out13_startofpacket (),                            // (terminated)
		.out13_endofpacket   (),                            // (terminated)
		.out13_empty         (),                            // (terminated)
		.out13_channel       (),                            // (terminated)
		.out13_error         (),                            // (terminated)
		.out13_data          (),                            // (terminated)
		.out14_ready         (1'b1),                        // (terminated)
		.out14_valid         (),                            // (terminated)
		.out14_startofpacket (),                            // (terminated)
		.out14_endofpacket   (),                            // (terminated)
		.out14_empty         (),                            // (terminated)
		.out14_channel       (),                            // (terminated)
		.out14_error         (),                            // (terminated)
		.out14_data          (),                            // (terminated)
		.out15_ready         (1'b1),                        // (terminated)
		.out15_valid         (),                            // (terminated)
		.out15_startofpacket (),                            // (terminated)
		.out15_endofpacket   (),                            // (terminated)
		.out15_empty         (),                            // (terminated)
		.out15_channel       (),                            // (terminated)
		.out15_error         (),                            // (terminated)
		.out15_data          ()                             // (terminated)
	);

	lab_PD1_sys_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                  (clk_clk),                                   //                                clk_clk.clk
		.my_masterB_reset_reset_bridge_in_reset_reset (~reset_reset_n),                            // my_masterB_reset_reset_bridge_in_reset.reset
		.my_masterB_m0_address                        (my_masterb_m0_address),                     //                          my_masterB_m0.address
		.my_masterB_m0_waitrequest                    (my_masterb_m0_waitrequest),                 //                                       .waitrequest
		.my_masterB_m0_write                          (my_masterb_m0_write),                       //                                       .write
		.my_masterB_m0_writedata                      (my_masterb_m0_writedata),                   //                                       .writedata
		.ST_ALU_0_s0_write                            (mm_interconnect_0_st_alu_0_s0_write),       //                            ST_ALU_0_s0.write
		.ST_ALU_0_s0_writedata                        (mm_interconnect_0_st_alu_0_s0_writedata),   //                                       .writedata
		.ST_ALU_0_s0_waitrequest                      (mm_interconnect_0_st_alu_0_s0_waitrequest), //                                       .waitrequest
		.ST_ALU_1_s0_write                            (mm_interconnect_0_st_alu_1_s0_write),       //                            ST_ALU_1_s0.write
		.ST_ALU_1_s0_writedata                        (mm_interconnect_0_st_alu_1_s0_writedata),   //                                       .writedata
		.ST_ALU_1_s0_waitrequest                      (mm_interconnect_0_st_alu_1_s0_waitrequest)  //                                       .waitrequest
	);

	lab_PD1_sys_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                                  (clk_clk),                                           //                                clk_clk.clk
		.my_masterA_reset_reset_bridge_in_reset_reset (~reset_reset_n),                                    // my_masterA_reset_reset_bridge_in_reset.reset
		.my_masterA_m0_address                        (my_mastera_m0_address),                             //                          my_masterA_m0.address
		.my_masterA_m0_waitrequest                    (my_mastera_m0_waitrequest),                         //                                       .waitrequest
		.my_masterA_m0_write                          (my_mastera_m0_write),                               //                                       .write
		.my_masterA_m0_writedata                      (my_mastera_m0_writedata),                           //                                       .writedata
		.MM_Stream_source_s0_write                    (mm_interconnect_1_mm_stream_source_s0_write),       //                    MM_Stream_source_s0.write
		.MM_Stream_source_s0_writedata                (mm_interconnect_1_mm_stream_source_s0_writedata),   //                                       .writedata
		.MM_Stream_source_s0_waitrequest              (mm_interconnect_1_mm_stream_source_s0_waitrequest)  //                                       .waitrequest
	);

	lab_PD1_sys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (0),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (0),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk   (clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset (~reset_reset_n),                // in_rst_0.reset
		.in_0_data      (st_splitter_out4_data),         //     in_0.data
		.in_0_valid     (st_splitter_out4_valid),        //         .valid
		.in_0_ready     (st_splitter_out4_ready),        //         .ready
		.out_0_data     (avalon_st_adapter_out_0_data),  //    out_0.data
		.out_0_valid    (avalon_st_adapter_out_0_valid)  //         .valid
	);

endmodule
