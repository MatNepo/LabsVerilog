
module lab_PD3_extra_task (
	clk_clk,
	reset_reset_n,
	dout_a_export,
	dout_b_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	dout_a_export;
	output	[31:0]	dout_b_export;
endmodule
