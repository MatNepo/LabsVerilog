
module Lab5_nios (
	clk_clk,
	led_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	led_export;
	input		reset_reset_n;
endmodule
