
module Lab1_task1_nios (
	clk_clk,
	led_export,
	reset_reset_n,
	sw_export);	

	input		clk_clk;
	output	[7:0]	led_export;
	input		reset_reset_n;
	input		sw_export;
endmodule
