// Sp_1.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Sp_1 (
		input  wire       source_clk, // source_clk.clk
		output wire [0:0] source      //    sources.source
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("SP 0"),
		.probe_width             (0),
		.source_width            (1),
		.source_initial_value    ("1"),
		.enable_metastability    ("YES")
	) in_system_sources_probes_0 (
		.source     (source),     //    sources.source
		.source_clk (source_clk), // source_clk.clk
		.source_ena (1'b1)        // (terminated)
	);

endmodule
